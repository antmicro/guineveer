// SPDX-License-Identifier: Apache-2.0
// Copyright (c) 2025-2026 Antmicro <www.antmicro.com>

`define HEX_FILE0 ""
`define HEX_FILE1 ""
