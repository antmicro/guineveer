`define HEX_FILE0 ""
`define HEX_FILE1 ""
